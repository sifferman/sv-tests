// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: arrays-packed-quering-functions-dimensions
:description: Test quering functions support on packed arrays
:tags: 7.11 7.4.1
:type: simulation elaboration parsing
*/
module top ();

bit [7:0] arr;

initial begin
	$svt_assert("(%d == 1)", $dimensions(arr));
end

endmodule
