// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: itor_function
:description: $itor test
:tags: 20.5
:type: simulation elaboration parsing
*/

module top();

initial begin
	$svt_assert("(%f == 20.0)", $itor(20));
end

endmodule
