// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: dyn-arr-basic
:description: Test dynamic arrays support
:tags: 7.5
:unsynthesizable: 1
*/
module top ();

bit [7:0] arr[];

endmodule
