// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: associative-arrays-integral
:description: Test associative arrays support
:tags: 7.8.4 7.8
:unsynthesizable: 1
*/
module top ();

int arr [ integer ];

endmodule
